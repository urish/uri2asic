magic
tech sky130A
timestamp 1638034600
<< nwell >>
rect -40 -195 205 -55
<< nmos >>
rect 40 0 55 65
<< pmos >>
rect 40 -140 55 -75
<< ndiff >>
rect 0 45 40 65
rect 0 25 5 45
rect 25 25 40 45
rect 0 0 40 25
rect 55 30 90 65
rect 55 10 65 30
rect 85 10 90 30
rect 55 0 90 10
<< pdiff >>
rect 0 -100 40 -75
rect 0 -120 5 -100
rect 25 -120 40 -100
rect 0 -140 40 -120
rect 55 -85 95 -75
rect 55 -105 70 -85
rect 90 -105 95 -85
rect 55 -140 95 -105
<< ndiffc >>
rect 5 25 25 45
rect 65 10 85 30
<< pdiffc >>
rect 5 -120 25 -100
rect 70 -105 90 -85
<< nsubdiff >>
rect 125 -145 180 -140
rect 125 -170 140 -145
rect 165 -170 180 -145
rect 125 -175 180 -170
<< nsubdiffcont >>
rect 140 -170 165 -145
<< poly >>
rect 40 65 55 90
rect 40 -15 55 0
rect 15 -25 55 -15
rect 15 -45 20 -25
rect 40 -45 55 -25
rect 15 -55 55 -45
rect 40 -75 55 -55
rect 40 -175 55 -140
<< polycont >>
rect 20 -45 40 -25
<< locali >>
rect -15 50 30 55
rect -55 45 30 50
rect -35 25 5 45
rect 25 25 30 45
rect -55 20 30 25
rect -15 10 30 20
rect 65 35 95 40
rect 65 30 115 35
rect 85 10 115 30
rect 65 0 115 10
rect 75 -15 115 0
rect -25 -25 55 -20
rect -5 -45 20 -25
rect 40 -45 55 -25
rect -25 -50 55 -45
rect 75 -40 95 -15
rect 75 -70 115 -40
rect 60 -85 115 -70
rect -15 -95 30 -90
rect -40 -100 30 -95
rect -20 -120 5 -100
rect 25 -120 30 -100
rect 60 -105 70 -85
rect 90 -105 115 -85
rect 60 -110 115 -105
rect 75 -120 115 -110
rect -40 -125 30 -120
rect -15 -140 30 -125
rect -15 -145 180 -140
rect -15 -170 140 -145
rect 165 -170 180 -145
rect -15 -175 180 -170
<< viali >>
rect -55 25 -35 45
rect -25 -45 -5 -25
rect 95 -40 115 -15
rect -40 -120 -20 -100
<< metal1 >>
rect -80 45 -25 50
rect -80 25 -55 45
rect -35 25 -25 45
rect -80 20 -25 25
rect 85 -15 160 -10
rect -50 -25 5 -20
rect -50 -45 -25 -25
rect -5 -45 5 -25
rect 85 -40 95 -15
rect 115 -40 160 -15
rect 85 -45 160 -40
rect -50 -50 5 -45
rect -80 -100 -10 -95
rect -80 -120 -40 -100
rect -20 -120 -10 -100
rect -80 -125 -10 -120
<< labels >>
rlabel metal1 120 -45 160 -10 1 Vout
rlabel metal1 -80 20 -55 50 1 Vss
rlabel metal1 -80 -125 -55 -95 1 Vdd
rlabel metal1 -50 -50 -25 -20 1 gate
<< end >>
