`default_nettype none
`timescale 1ns/1ps
module seven_segment (
    input wire          clk,
    input wire          reset,
    input wire          load,
    input wire [3:0]    ten_count,
    input wire [3:0]    unit_count,
    output reg [6:0]    segments,
    output reg          digit
);

reg [3:0]ten;
reg [3:0]unit;
wire [3:0]digit_value = digit ? ten : unit;

always @(*) begin
    case(digit_value)
        //                7654321
        0:  segments = 7'b0111111;
        1:  segments = 7'b0000110;
        2:  segments = 7'b1011011;
        3:  segments = 7'b1001111;
        4:  segments = 7'b1100110;
        5:  segments = 7'b1101101;
        6:  segments = 7'b1111100;
        7:  segments = 7'b0000111;
        8:  segments = 7'b1111111;
        9:  segments = 7'b1100111;
        default:    
            segments = 7'b0000000;
    endcase
end

always @(posedge clk) begin
    if (reset) begin
        ten <= 4'hf;
        unit <= 4'hf;
        digit <= 0;
    end else begin
        digit <= !digit;
        if (load) begin
            ten <= ten_count;
            unit <= unit_count;
        end
    end
end

endmodule
