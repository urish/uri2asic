.ends

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create a resistor between the MOSFET output and VGND
*R VPWR VOUT 10k

* create pulse
Vin GATE VGND pulse(0 1.8 1p 10p 10p 1n 2n)
.tran 10p 4n 0

.control
run
set color0 = white
set color1 = black
plot Vout GATE
.endc

.end
