MOSFET Simulation
* this file edited to remove everything not in tt lib
.lib "./sky130_fd_pr/models/sky130.lib.spice" tt

* instantiate the inverter
Xmosfet VPWR VGND GATE VOUT VGND X0

.subckt X0 Vdd Vss gate Vout VSUBS
* NGSPICE file created from mosfet.ext - technology: sky130A


* Top level circuit mosfet

X0 Vout gate Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Vout gate Vss VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
C0 Vdd Vss 0.04fF
C1 Vout Vss 0.03fF
C2 Vdd gate 0.12fF
C3 Vout gate 0.06fF
C4 Vss gate 0.09fF
C5 Vdd Vout 0.14fF
C6 Vout VSUBS 0.23fF
C7 Vss VSUBS 0.15fF
C8 gate VSUBS 0.27fF
C9 Vdd VSUBS 0.74fF


.ends

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create a resistor between the MOSFET output and VGND
*R VPWR VOUT 10k

* create pulse
Vin GATE VGND pulse(0 1.8 1p 10p 10p 1n 2n)
.tran 10p 4n 0

.control
run
set color0 = white
set color1 = black
plot Vout GATE
.endc

.end
